../../sva/rf_stage.sv