../../sva/eth_top.sv