../../sva/mips_dvc.sv