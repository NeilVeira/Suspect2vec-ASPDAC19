../../sva/ctl_fsm.sv