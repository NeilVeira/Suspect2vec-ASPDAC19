../../sva/VennsaChecker.sv