../../sva/spi_top.sv