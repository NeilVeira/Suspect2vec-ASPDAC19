../../sva/vga_fifo.sv