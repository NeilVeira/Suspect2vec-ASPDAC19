../../sva/vga_top.sv