../../sva/vga_colproc.sv