../../sva/wb_master.sv