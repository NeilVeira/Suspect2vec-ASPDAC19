../../sva/mips_sys.sv