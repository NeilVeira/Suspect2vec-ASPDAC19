../../sva/check.sv