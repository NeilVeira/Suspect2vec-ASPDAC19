../../sva/vga_pgen.sv