../../sva/fifo4.sv