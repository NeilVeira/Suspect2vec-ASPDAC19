../../sva/exec_stage.sv