../../sva/wb_slave.sv